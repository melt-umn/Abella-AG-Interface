grammar interface_:toAbella;

imports interface_:common:abstractSyntax;

exports interface_:toAbella:concreteSyntax;
exports interface_:toAbella:abstractSyntax;