grammar toAbella;

exports toAbella:concreteSyntax;
exports toAbella:abstractSyntax;