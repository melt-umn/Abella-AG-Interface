grammar interface_:fromAbella:abstractSyntax;

