grammar interface_:common;

exports interface_:common:concreteSyntax;
exports interface_:common:abstractSyntax;

