grammar interface_:thm_interface_file;


exports interface_:thm_interface_file:concreteSyntax;
exports interface_:thm_interface_file:abstractSyntax;

