grammar interface_:toAbella:abstractSyntax;


attribute
   cleanUpCommands, numCleanUpCommands,
   nextStateIn, nextStateOut,
   treeTys
occurs on ProofState;


aspect production proofInProgress
top::ProofState ::=
   subgoalNum::[Integer] currGoal::CurrentGoal futureGoals::[Subgoal]
{
  --Clean up attribute accesses to be equal
  --(hyp name, tree name, attr name, type name, value of attr)
  local attrAccessHyps::[(String, String, String, String, Term)] =
        foldr(
          \ p::(String, Metaterm)
            rest::[(String, String, String, String, Term)] ->
            case p.1, decorate p.2 with {silverContext = top.silverContext;} of
            | hyp,
              termMetaterm(applicationTerm(nameTerm(access, _),
                             consTermList(nameTerm(treeName, _),
                             consTermList(nameTerm(treeNode, _),
                             singleTermList(val)))), _)
              when isAccessRelation(access) ->
              (hyp, treeName,
               accessRelationToAttr(access),
               accessRelationToType(access), new(val))::rest
            | _, _ -> rest
            end,
          [], currGoal.hypList);
  local sortedAttrAccessHyps::[(String, String, String, String, Term)] =
        sortBy(\ p1::(String, String, String, String, Term)
                 p2::(String, String, String, String, Term) ->
                 p1.3 < p2.3 || (p1.3 == p2.3 && p1.2 <= p2.2),
               attrAccessHyps);
  local groupedAttrAccesses::[[(String, String, String, String, Term)]] =
        groupBy(\ p1::(String, String, String, String, Term)
                  p2::(String, String, String, String, Term) ->
                  p1.2 == p2.2 && p1.3 == p2.3,
                sortedAttrAccessHyps);
  local cleanedAttrAccessGroups::[[(String, String, String, String, Term)]] =
        map(\ l::[(String, String, String, String, Term)] ->
              nubBy(\ p1::(String, String, String, String, Term)
                      p2::(String, String, String, String, Term) ->
                    p1.5.pp == p2.5.pp, l), groupedAttrAccesses);
  local cleanedAttrAccesses::[[(String, String, String, String, Term)]] =
        filter(\ l::[(String, String, String, String, Term)] ->
                 length(l) > 1, cleanedAttrAccessGroups);
  --We can only do one clean up at a time, since each one might
  --   eliminate the goal based on impossibility
  --We can do the rest later, if we don't remove the goal
  local attrAccessCmd::String =
        case head(cleanedAttrAccesses) of
        | (hyp1, _, attr, ty, _)::(hyp2, _, _, _, _)::_ ->
          applyTactic(noHint(), nothing(),
                      clearable(false, accessUniqueThm(attr, ty), []),
                      [hypApplyArg(hyp1, []),
                       hypApplyArg(hyp2, [])], []).pp
        | _ -> error("Impossible after filtration")
        end;

  --Clean up local attribute accesses to be equal
  --(hyp name, tree name, prod name, attr name, type name, value of attr)
  local localAccessHyps::[(String, String, String, String, String, Term)] =
        foldr(
          \ p::(String, Metaterm)
            rest::[(String, String, String, String, String, Term)] ->
            case p.1, decorate p.2 with {silverContext = top.silverContext;} of
            | hyp,
              termMetaterm(applicationTerm(nameTerm(access, _),
                             consTermList(nameTerm(treeName, _),
                             consTermList(nameTerm(treeNode, _),
                             singleTermList(val)))), _)
              when isLocalAccessRelation(access) ->
              (hyp, treeName,
               localAccessToProd(access),
               localAccessToAttr(access),
               localAccessToType(access).pp, new(val))::rest
            | _, _ -> rest
            end,
          [], currGoal.hypList);
  local sortedLocalAccessHyps::[(String, String, String, String, String, Term)] =
        sortBy(\ p1::(String, String, String, String, String, Term)
                 p2::(String, String, String, String, String, Term) ->
                 p1.4 < p2.4 || (p1.4 == p2.4 && p1.2 <= p2.2),
               localAccessHyps);
  local groupedLocalAccesses::[[(String, String, String, String, String, Term)]] =
        groupBy(\ p1::(String, String, String, String, String, Term)
                  p2::(String, String, String, String, String, Term) ->
                  p1.2 == p2.2 && p1.3 == p2.3 && p1.4 == p2.4,
                sortedLocalAccessHyps);
  local cleanedLocalAccessGroups::[[(String, String, String, String, String, Term)]] =
        map(\ l::[(String, String, String, String, String, Term)] ->
              nubBy(\ p1::(String, String, String, String, String, Term)
                      p2::(String, String, String, String, String, Term) ->
                    p1.6.pp == p2.6.pp, l), groupedLocalAccesses);
  local cleanedLocalAccesses::[[(String, String, String, String, String, Term)]] =
        filter(\ l::[(String, String, String, String, String, Term)] ->
                 length(l) > 1, cleanedLocalAccessGroups);
  --We can only do one clean up at a time, since each one might
  --   eliminate the goal based on impossibility
  --We can do the rest later, if we don't remove the goal
  local localAccessCmd::String =
        case head(cleanedLocalAccesses) of
        | (hyp1, _, prod, attr, ty, _)::(hyp2, _, _, _, _, _)::_ ->
          applyTactic(noHint(), nothing(),
                      clearable(false, localAccessUniqueThm(prod, attr, ty), []),
                      [hypApplyArg(hyp1, []),
                       hypApplyArg(hyp2, [])], []).pp
        | _ -> error("Impossible after filtration")
        end;

  --Clean up cases with impossible tree forms which come from equations
  --   for local attributes
  --We need to hide these cases to hide the encoding of the AG
  --(exists <Children>, <prod>(<Children'>) = <prod>(<Children>)) -> false
  local impossibleEqHyps::[String] =
        foldr(\ p::(String, Metaterm) rest::[String] ->
                case p.1, decorate p.2 with {silverContext = top.silverContext;} of
                --TODO need to handle non-tree children
                | hyp,
                  impliesMetaterm(
                     bindingMetaterm(
                        existsBinder(),
                        children,
                        eqMetaterm(
                           applicationTerm(nameTerm(prod1, _), args1),
                           applicationTerm(nameTerm(prod2, _), args2))),
                     falseMetaterm())
                  when isProd(prod1) && prod1 == prod2 ->
                  hyp::rest
                | hyp,
                  impliesMetaterm(
                     bindingMetaterm(
                        existsBinder(),
                        children,
                        eqMetaterm(
                           nameTerm(prod1, _),
                           nameTerm(prod2, _))),
                     falseMetaterm())
                  when isProd(prod1) && prod1 == prod2 -> hyp::rest
                | _, _ -> rest
                end,
              [], currGoal.hypList);
  local impossibleEqHypsCmd::String =
        let name::String = "$F_" ++ toString(genInt())
        in
          name ++ ": assert false.  " ++
          "backchain " ++ head(impossibleEqHyps) ++ ".  " ++
          "case " ++ name ++ ".  "
        end;

  top.cleanUpCommands =
      if null(cleanedAttrAccesses)
      then if null(cleanedLocalAccesses)
           then if null(impossibleEqHyps)
                then ""
                else impossibleEqHypsCmd
           else localAccessCmd
      else attrAccessCmd;
  top.numCleanUpCommands =
      if null(cleanedAttrAccesses)
      then if null(cleanedLocalAccesses)
           then if null(impossibleEqHyps)
                then 0
                else 3
           else 1
      else 1;

  top.nextStateOut = top.nextStateIn;
  currGoal.knownDecoratedTrees = top.gatheredDecoratedTrees;
}


aspect production noProof
top::ProofState ::=
{
  top.cleanUpCommands = "";
  top.numCleanUpCommands = 0;

  top.nextStateOut = top.nextStateIn;
}


aspect production extensible_proofInProgress
top::ProofState ::=
     currentProofState::ProofState
     originalTheorems::[(String, Metaterm)]
     numProds::[(String, Integer)]
{
  --names for the split theorems
  local newThmNames::[String] =
        flatMap(\ p::(String, Integer) ->
           map(\ i::Integer -> "$" ++ colonsToEncoded(p.1) ++ "_$_" ++ toString(i),
               range(1, p.2 + 1)),
           numProds);
  local isDone::Boolean =
        case currentProofState of
        | proofInProgress(_, _, _) -> false
        | proofCompleted() -> true
        | proofAborted() -> true
        | noProof() ->
          error("Should not have extensible_proofInProgress of noProof")
        end;
  local shouldDeclare::Boolean =
        case currentProofState of
        | proofInProgress(_, _, _) -> false
        | proofCompleted() -> true
        | proofAborted() -> false
        | noProof() ->
          error("Should not have extensible_proofInProgress of noProof")
        end;
  top.cleanUpCommands =
      if isDone && shouldDeclare
      then --split, declare, and skip.
           splitTheorem(
              extensible_theorem_name(colonsToEncoded(head(originalTheorems).1),
                 top.silverContext.currentGrammar),
              newThmNames).pp ++
           foldr(\ p::(String, Metaterm) rest::String ->
                   theoremDeclaration(colonsToEncoded(p.1), [], p.2).pp ++ "  " ++
                   skipTactic().pp ++ "\n" ++ rest,
                 "", originalTheorems)
      else currentProofState.cleanUpCommands;
  top.numCleanUpCommands =
      if isDone && shouldDeclare
      then 1 + 2 * length(originalTheorems)
      else currentProofState.numCleanUpCommands;

  top.nextStateOut =
      if isDone
      then top.nextStateIn
      else extensible_proofInProgress(
              top.nextStateIn, originalTheorems, numProds);}


abstract production obligation_proofInProgress
top::ProofState ::=
     currentProofState::ProofState
     originalTheorems::[(String, Metaterm)]
     numProds::[(String, Integer)]
{
  local isDone::Boolean =
        case currentProofState of
        | proofInProgress(_, _, _) -> false
        | proofCompleted() -> true
        | proofAborted() -> true
        | noProof() ->
          error("Should not have obligation_proofInProgress of noProof")
        end;
  local shouldDeclare::Boolean =
        case currentProofState of
        | proofInProgress(_, _, _) -> false
        | proofCompleted() -> true
        | proofAborted() -> false
        | noProof() ->
          error("Should not have obligation_proofInProgress of noProof")
        end;
  top.nextStateOut =
      if isDone
      then top.nextStateIn
      else obligation_proofInProgress(
              top.nextStateIn, originalTheorems, numProds);

  forwards to extensible_proofInProgress(currentProofState,
                 originalTheorems, numProds);
}



attribute
   knownDecoratedTrees,
   treeTys
occurs on CurrentGoal;

aspect production currentGoal
top::CurrentGoal ::= vars::[String] ctx::Context goal::Metaterm
{

}



attribute
   knownDecoratedTrees,
   treeTys
occurs on Context;

aspect production emptyContext
top::Context ::=
{
  
}


aspect production singleContext
top::Context ::= h::Hypothesis
{
  
}


aspect production branchContext
top::Context ::= c1::Context c2::Context
{
  
}



attribute
   knownDecoratedTrees,
   treeTys
occurs on Hypothesis;

aspect production metatermHyp
top::Hypothesis ::= name::String body::Metaterm
{
  
}

