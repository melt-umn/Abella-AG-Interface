grammar interface_:fromAbella;

imports interface_:common;

exports interface_:fromAbella:concreteSyntax;
exports interface_:fromAbella:abstractSyntax;