grammar fromAbella;

exports fromAbella:concreteSyntax;
exports fromAbella:abstractSyntax;