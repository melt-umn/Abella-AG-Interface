grammar interface_:thmInterfaceFile;


exports interface_:thmInterfaceFile:concreteSyntax;
exports interface_:thmInterfaceFile:abstractSyntax;

