grammar interface_:toAbella;

imports interface_:common;

exports interface_:toAbella:concreteSyntax;
exports interface_:toAbella:abstractSyntax;