grammar toAbella:abstractSyntax;


synthesized attribute pp::String;

